module sum( 
input [15:0] a, 
input [15:0] b, 
output [15:0] res 
); 

assign res = a + b; 

endmodule
